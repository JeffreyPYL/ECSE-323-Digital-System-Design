library verilog;
use verilog.vl_types.all;
entity g19_Envelope_vlg_vec_tst is
end g19_Envelope_vlg_vec_tst;
